   output                     bootrom_r_en,
   output [`BOOTROM_ADDR_W-2-1:0]       bootrom_addr,
   input [`DATA_W-1:0]        bootrom_r_data,

