   output                     bootrom_r_en,
   output [`ADDR_W-1:0]       bootrom_addr,
   input [`DATA_W-1:0]        bootrom_r_data,

