        .bootrom_r_en(bootrom_r_en),
        .bootrom_addr(bootrom_addr),
        .bootrom_r_data(bootrom_r_data),
        
