`timescale 1ns / 1ps
`include "system.vh"
`include "axi.vh"

module top_system(
	          input         c0_sys_clk_clk_p, 
                  input         c0_sys_clk_clk_n, 
	          input         reset,

	          //uart
	          output        uart_txd,
	          input         uart_rxd,

`ifdef USE_DDR
                  output        c0_ddr4_act_n,
                  output [16:0] c0_ddr4_adr,
                  output [1:0]  c0_ddr4_ba,
                  output [0:0]  c0_ddr4_bg,
                  output [0:0]  c0_ddr4_cke,
                  output [0:0]  c0_ddr4_odt,
                  output [0:0]  c0_ddr4_cs_n,
                  output [0:0]  c0_ddr4_ck_t,
                  output [0:0]  c0_ddr4_ck_c,
                  output        c0_ddr4_reset_n,
                  inout [3:0]   c0_ddr4_dm_dbi_n,
                  inout [31:0]  c0_ddr4_dq,
                  inout [3:0]   c0_ddr4_dqs_c,
                  inout [3:0]   c0_ddr4_dqs_t, 
`endif                  
		  output        trap
		  );

`ifdef USE_DDR
   //
   // AXI INTERCONNECT
   //
                         
   // SYSTEM/SLAVE SIDE
   // address write
   wire [2*1-1:0]           sys_axi_awid;
   wire [2*`DDR_ADDR_W-1:0] sys_axi_awaddr;
   wire [2*8-1:0]           sys_axi_awlen;
   wire [2*3-1:0]           sys_axi_awsize;
   wire [2*2-1:0]           sys_axi_awburst;
   wire [2*1-1:0]           sys_axi_awlock;
   wire [2*4-1:0]           sys_axi_awcache;
   wire [2*3-1:0]           sys_axi_awprot;
   wire [2*4-1:0]           sys_axi_awqos;
   wire [2*1-1:0]           sys_axi_awvalid;
   wire [2*1-1:0]           sys_axi_awready;
   //write
   wire [2*32-1:0]          sys_axi_wdata;
   wire [2*4-1:0]           sys_axi_wstrb;
   wire [2*1-1:0]           sys_axi_wlast;
   wire [2*1-1:0]           sys_axi_wvalid;
   wire [2*1-1:0]           sys_axi_wready;
   //write response
   wire [2*1-1:0]           sys_axi_bid;
   wire [2*2-1:0]           sys_axi_bresp;
   wire [2*1-1:0]           sys_axi_bvalid;
   wire [2*1-1:0]           sys_axi_bready;
   //address read
   wire [2*1-1:0]           sys_axi_arid;
   wire [2*`DDR_ADDR_W-1:0] sys_axi_araddr;
   wire [2*8-1:0]           sys_axi_arlen;
   wire [2*3-1:0]           sys_axi_arsize;
   wire [2*2-1:0]           sys_axi_arburst;
   wire [2*1-1:0]           sys_axi_arlock;
   wire [2*4-1:0]           sys_axi_arcache;
   wire [2*3-1:0]           sys_axi_arprot;
   wire [2*4-1:0]           sys_axi_arqos;
   wire [2*1-1:0]           sys_axi_arvalid;
   wire [2*1-1:0]           sys_axi_arready;
   //read
   wire [2*1-1:0]           sys_axi_rid;
   wire [2*`DATA_W-1:0]     sys_axi_rdata;   
   wire [2*2-1:0]           sys_axi_rresp;   
   wire [2*1-1:0]           sys_axi_rlast;
   wire [2*1-1:0]           sys_axi_rvalid;
   wire [2*1-1:0]           sys_axi_rready;

   // DDR/MASTER SIDE
   `AXI4_IF_WIRE(ddr)
`endif


   //
   // CLOCK MANAGEMENT
   //

   //system clock
   wire 			sys_clk;
   
`ifdef USE_DDR
   wire                         ddr_aclk;
`else 
   clock_wizard #(
		  .OUTPUT_PER(10),
		  .INPUT_PER(4)
		  )
   clk_250_to_100_MHz(
		      .clk_in1_p(c0_sys_clk_clk_p),
		      .clk_in1_n(c0_sys_clk_clk_n),
		      .clk_out1(sys_clk)
		      );
`endif
   
   //ddr clock output from ddr ctrl 
 


   //   
   // RESET MANAGEMENT
   //

   //system reset
 
   wire                         sys_rst;

`ifdef USE_DDR
   wire                         init_calib_complete;
   wire                         sys_rstn;

   assign sys_rst  = ~sys_rstn;
`else
   reg [15:0] 			rst_cnt;
   reg                          sys_rst_int;
   
   always @(posedge sys_clk, posedge reset)
     if(reset) begin
        sys_rst_int <= 1'b0;
        rst_cnt <= 16'hFFFF;
     end else begin 
        if(rst_cnt != 16'h0)
          rst_cnt <= rst_cnt - 1'b1;
        sys_rst_int <= (rst_cnt != 16'h0);
     end

   assign sys_rst = sys_rst_int;
   
`endif

`ifdef USE_DDR
   //AXI DDR side reset (ddr_arst) : generated by MIG itself
   wire                         ddr_arstn;   
   wire                         ddr_ui_clk;
`endif
   

   //
   // DDR CONTROLLER
   //
                 
`ifdef USE_DDR   
   ddr4_0 ddr4_ram 
     (
      .sys_rst                (reset),
      .c0_sys_clk_p           (c0_sys_clk_clk_p),
      .c0_sys_clk_n           (c0_sys_clk_clk_n),

      .dbg_clk                (),
      .dbg_bus                (),
      
      //EXTERNAL SIDE
      .c0_ddr4_act_n          (c0_ddr4_act_n),
      .c0_ddr4_adr            (c0_ddr4_adr),
      .c0_ddr4_ba             (c0_ddr4_ba),
      .c0_ddr4_bg             (c0_ddr4_bg),
      .c0_ddr4_cke            (c0_ddr4_cke),
      .c0_ddr4_odt            (c0_ddr4_odt),
      .c0_ddr4_cs_n           (c0_ddr4_cs_n),
      .c0_ddr4_ck_t           (c0_ddr4_ck_t),
      .c0_ddr4_ck_c           (c0_ddr4_ck_c),
      .c0_ddr4_reset_n        (c0_ddr4_reset_n),
      .c0_ddr4_dm_dbi_n       (c0_ddr4_dm_dbi_n),
      .c0_ddr4_dq             (c0_ddr4_dq),
      .c0_ddr4_dqs_c          (c0_ddr4_dqs_c),
      .c0_ddr4_dqs_t          (c0_ddr4_dqs_t),
      .c0_init_calib_complete (init_calib_complete),
      
      //generated clocks and resets
      .c0_ddr4_ui_clk         (ddr_ui_clk),
      .c0_ddr4_ui_clk_sync_rst(ddr_ui_rst),
      .addn_ui_clkout1        (sys_clk),

      //USER AXI INTERFACE
      .c0_ddr4_aresetn        (ddr_arstn),

      `AXI4_IF_PORTMAP(c0_ddr4_s_,ddr_)
      );   


   axi_interconnect_0 cache2ddr 
     (
      .INTERCONNECT_ACLK     (ddr_ui_clk),
      .INTERCONNECT_ARESETN  (~(ddr_ui_rst | ~init_calib_complete)),
      
      //
      // SYSTEM SIDE
      //
      .S00_AXI_ARESET_OUT_N (sys_rstn),
      .S00_AXI_ACLK         (sys_clk),
      
     //Write address
      .S00_AXI_AWID         (sys_axi_awid[0*1+:1]),
      .S00_AXI_AWADDR       (sys_axi_awaddr[0*`DDR_ADDR_W+:`DDR_ADDR_W]),
      .S00_AXI_AWLEN        (sys_axi_awlen[0*8+:8]),
      .S00_AXI_AWSIZE       (sys_axi_awsize[0*3+:3]),
      .S00_AXI_AWBURST      (sys_axi_awburst[0*2+:2]),
      .S00_AXI_AWLOCK       (sys_axi_awlock[0*1+:1]),
      .S00_AXI_AWCACHE      (sys_axi_awcache[0*4+:4]),
      .S00_AXI_AWPROT       (sys_axi_awprot[0*3+:3]),
      .S00_AXI_AWQOS        (sys_axi_awqos[0*4+:4]),
      .S00_AXI_AWVALID      (sys_axi_awvalid[0*1+:1]),
      .S00_AXI_AWREADY      (sys_axi_awready[0*1+:1]),

      //Write data
      .S00_AXI_WDATA        (sys_axi_wdata[0*32+:32]),
      .S00_AXI_WSTRB        (sys_axi_wstrb[0*4+:4]),
      .S00_AXI_WLAST        (sys_axi_wlast[0*1+:1]),
      .S00_AXI_WVALID       (sys_axi_wvalid[0*1+:1]),
      .S00_AXI_WREADY       (sys_axi_wready[0*1+:1]),
      
      //Write response
      .S00_AXI_BID           (sys_axi_bid[0*1+:1]),
      .S00_AXI_BRESP         (sys_axi_bresp[0*2+:2]),
      .S00_AXI_BVALID        (sys_axi_bvalid[0*1+:1]),
      .S00_AXI_BREADY        (sys_axi_bready[0*1+:1]),
      
      //Read address
      .S00_AXI_ARID         (sys_axi_arid[0*1+:1]),
      .S00_AXI_ARADDR       (sys_axi_araddr[0*`DDR_ADDR_W+:`DDR_ADDR_W]),
      .S00_AXI_ARLEN        (sys_axi_arlen[0*8+:8]),
      .S00_AXI_ARSIZE       (sys_axi_arsize[0*3+:3]),
      .S00_AXI_ARBURST      (sys_axi_arburst[0*2+:2]),
      .S00_AXI_ARLOCK       (sys_axi_arlock[0*1+:1]),
      .S00_AXI_ARCACHE      (sys_axi_arcache[0*4+:4]),
      .S00_AXI_ARPROT       (sys_axi_arprot[0*3+:3]),
      .S00_AXI_ARQOS        (sys_axi_arqos[0*4+:4]),
      .S00_AXI_ARVALID      (sys_axi_arvalid[0*1+:1]),
      .S00_AXI_ARREADY      (sys_axi_arready[0*1+:1]),
      
      //Read data
      .S00_AXI_RID          (sys_axi_rid[0*1+:1]),
      .S00_AXI_RDATA        (sys_axi_rdata[0*`DATA_W+:`DATA_W]),
      .S00_AXI_RRESP        (sys_axi_rresp[0*2+:2]),
      .S00_AXI_RLAST        (sys_axi_rlast[0*1+:1]),
      .S00_AXI_RVALID       (sys_axi_rvalid[0*1+:1]),
      .S00_AXI_RREADY       (sys_axi_rready[0*1+:1]),

      .S01_AXI_ARESET_OUT_N (),
      .S01_AXI_ACLK         (sys_clk),
      
      //Write address
      .S01_AXI_AWID         (sys_axi_awid[1*1+:1]),
      .S01_AXI_AWADDR       (sys_axi_awaddr[1*`DDR_ADDR_W+:`DDR_ADDR_W]),
      .S01_AXI_AWLEN        (sys_axi_awlen[1*8+:8]),
      .S01_AXI_AWSIZE       (sys_axi_awsize[1*3+:3]),
      .S01_AXI_AWBURST      (sys_axi_awburst[1*2+:2]),
      .S01_AXI_AWLOCK       (sys_axi_awlock[1*1+:1]),
      .S01_AXI_AWCACHE      (sys_axi_awcache[1*4+:4]),
      .S01_AXI_AWPROT       (sys_axi_awprot[1*3+:3]),
      .S01_AXI_AWQOS        (sys_axi_awqos[1*4+:4]),
      .S01_AXI_AWVALID      (sys_axi_awvalid[1*1+:1]),
      .S01_AXI_AWREADY      (sys_axi_awready[1*1+:1]),

      //Write data
      .S01_AXI_WDATA        (sys_axi_wdata[1*32+:32]),
      .S01_AXI_WSTRB        (sys_axi_wstrb[1*4+:4]),
      .S01_AXI_WLAST        (sys_axi_wlast[1*1+:1]),
      .S01_AXI_WVALID       (sys_axi_wvalid[1*1+:1]),
      .S01_AXI_WREADY       (sys_axi_wready[1*1+:1]),
      
      //Write response
      .S01_AXI_BID           (sys_axi_bid[1*1+:1]),
      .S01_AXI_BRESP         (sys_axi_bresp[1*2+:2]),
      .S01_AXI_BVALID        (sys_axi_bvalid[1*1+:1]),
      .S01_AXI_BREADY        (sys_axi_bready[1*1+:1]),
      
      //Read address
      .S01_AXI_ARID         (sys_axi_arid[1*1+:1]),
      .S01_AXI_ARADDR       (sys_axi_araddr[1*`DDR_ADDR_W+:`DDR_ADDR_W]),
      .S01_AXI_ARLEN        (sys_axi_arlen[1*8+:8]),
      .S01_AXI_ARSIZE       (sys_axi_arsize[1*3+:3]),
      .S01_AXI_ARBURST      (sys_axi_arburst[1*2+:2]),
      .S01_AXI_ARLOCK       (sys_axi_arlock[1*1+:1]),
      .S01_AXI_ARCACHE      (sys_axi_arcache[1*4+:4]),
      .S01_AXI_ARPROT       (sys_axi_arprot[1*3+:3]),
      .S01_AXI_ARQOS        (sys_axi_arqos[1*4+:4]),
      .S01_AXI_ARVALID      (sys_axi_arvalid[1*1+:1]),
      .S01_AXI_ARREADY      (sys_axi_arready[1*1+:1]),
      
      //Read data
      .S01_AXI_RID          (sys_axi_rid[1*1+:1]),
      .S01_AXI_RDATA        (sys_axi_rdata[1*`DATA_W+:`DATA_W]),
      .S01_AXI_RRESP        (sys_axi_rresp[1*2+:2]),
      .S01_AXI_RLAST        (sys_axi_rlast[1*1+:1]),
      .S01_AXI_RVALID       (sys_axi_rvalid[1*1+:1]),
      .S01_AXI_RREADY       (sys_axi_rready[1*1+:1]),
      //
      // DDR SIDE
      //

      .M00_AXI_ARESET_OUT_N  (ddr_arstn),
      .M00_AXI_ACLK          (ddr_ui_clk),
      
      //Write address
      .M00_AXI_AWID          (ddr_axi_awid),
      .M00_AXI_AWADDR        (ddr_axi_awaddr),
      .M00_AXI_AWLEN         (ddr_axi_awlen),
      .M00_AXI_AWSIZE        (ddr_axi_awsize),
      .M00_AXI_AWBURST       (ddr_axi_awburst),
      .M00_AXI_AWLOCK        (ddr_axi_awlock),
      .M00_AXI_AWCACHE       (ddr_axi_awcache),
      .M00_AXI_AWPROT        (ddr_axi_awprot),
      .M00_AXI_AWQOS         (ddr_axi_awqos),
      .M00_AXI_AWVALID       (ddr_axi_awvalid),
      .M00_AXI_AWREADY       (ddr_axi_awready),
      
      //Write data
      .M00_AXI_WDATA         (ddr_axi_wdata),
      .M00_AXI_WSTRB         (ddr_axi_wstrb),
      .M00_AXI_WLAST         (ddr_axi_wlast),
      .M00_AXI_WVALID        (ddr_axi_wvalid),
      .M00_AXI_WREADY        (ddr_axi_wready),
      
      //Write response
      .M00_AXI_BID           (ddr_axi_bid),
      .M00_AXI_BRESP         (ddr_axi_bresp),
      .M00_AXI_BVALID        (ddr_axi_bvalid),
      .M00_AXI_BREADY        (ddr_axi_bready),
      
      //Read address
      .M00_AXI_ARID         (ddr_axi_arid),
      .M00_AXI_ARADDR       (ddr_axi_araddr),
      .M00_AXI_ARLEN        (ddr_axi_arlen),
      .M00_AXI_ARSIZE       (ddr_axi_arsize),
      .M00_AXI_ARBURST      (ddr_axi_arburst),
      .M00_AXI_ARLOCK       (ddr_axi_arlock),
      .M00_AXI_ARCACHE      (ddr_axi_arcache),
      .M00_AXI_ARPROT       (ddr_axi_arprot),
      .M00_AXI_ARQOS        (ddr_axi_arqos),
      .M00_AXI_ARVALID      (ddr_axi_arvalid),
      .M00_AXI_ARREADY      (ddr_axi_arready),
      
      //Read data
      .M00_AXI_RID          (ddr_axi_rid),
      .M00_AXI_RDATA        (ddr_axi_rdata),
      .M00_AXI_RRESP        (ddr_axi_rresp),
      .M00_AXI_RLAST        (ddr_axi_rlast),
      .M00_AXI_RVALID       (ddr_axi_rvalid),
      .M00_AXI_RREADY       (ddr_axi_rready)
      );
`endif

   //
   // SYSTEM
   //
   system system 
     (
      .clk           (sys_clk),
      .reset         (sys_rst),
      .trap          (trap),

`ifdef USE_DDR
      `AXI4_IF_PORTMAP(m_,sys_),
`endif
      
      //UART
      .uart_txd      (uart_txd),
      .uart_rxd      (uart_rxd),
      .uart_rts      (),
      .uart_cts      (1'b1)
      );
   
endmodule
