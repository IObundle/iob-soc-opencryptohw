    // sram data ports
    .sram_enA   (sram_enA),
    .sram_addrA (sram_addrA),
    .sram_weA   (sram_weA),
    .sram_dinA  (sram_dinA),
    .sram_doutA (sram_doutA),

    // sram instruction ports
    .sram_enB   (sram_enB),
    .sram_addrB (sram_addrB),
    .sram_weB   (sram_weB),
    .sram_dinB  (sram_dinB),
    .sram_doutB (sram_doutB),
