`timescale 1ns / 1ps
`include "axi.vh"
`include "xversat.vh"
`include "xdefs.vh"

module M #(
      parameter ADDR_W = `ADDR_W,
      parameter DATA_W = `DATA_W,
      parameter AXI_ADDR_W = `AXI_ADDR_W
   )
   (

   input run,
   output done,

   input [DATA_W-1:0]              in0,
   input [DATA_W-1:0]              in1,
   input [DATA_W-1:0]              in2,
   input [DATA_W-1:0]              in3,
   input [DATA_W-1:0]              in4,
   input [DATA_W-1:0]              in5,
   input [DATA_W-1:0]              in6,
   input [DATA_W-1:0]              in7,
   input [DATA_W-1:0]              in8,
   input [DATA_W-1:0]              in9,
   input [DATA_W-1:0]              in10,
   input [DATA_W-1:0]              in11,
   input [DATA_W-1:0]              in12,
   input [DATA_W-1:0]              in13,
   input [DATA_W-1:0]              in14,
   input [DATA_W-1:0]              in15,
   output [DATA_W-1:0]             out0,
   output [DATA_W-1:0]             out1,
   output [DATA_W-1:0]             out2,
   output [DATA_W-1:0]             out3,
   output [DATA_W-1:0]             out4,
   output [DATA_W-1:0]             out5,
   output [DATA_W-1:0]             out6,
   output [DATA_W-1:0]             out7,
   output [DATA_W-1:0]             out8,
   output [DATA_W-1:0]             out9,
   output [DATA_W-1:0]             out10,
   output [DATA_W-1:0]             out11,
   output [DATA_W-1:0]             out12,
   output [DATA_W-1:0]             out13,
   output [DATA_W-1:0]             out14,
   output [DATA_W-1:0]             out15,
   input [31:0]     constant_0,
   input [31:0]     constant_1,
   input [31:0]     constant_2,
   input [31:0]     constant_3,
   input [31:0]     constant_4,
   input [31:0]     constant_5,
   input [31:0]     constant_6,
   input [31:0]     constant_7,
   input [31:0]     constant_8,
   input [31:0]     constant_9,
   input [31:0]     constant_10,
   input [31:0]     constant_11,
   input [31:0]     constant_12,
   input [31:0]     constant_13,
   input [31:0]     constant_14,
   input [31:0]     constant_15,
   input [31:0]     constant_16,
   input [31:0]     constant_17,
   input [31:0]     constant_18,
   input [31:0]     constant_19,
   input [31:0]     constant_20,
   input [31:0]     constant_21,
   input [31:0]     constant_22,
   input [31:0]     constant_23,
   input [31:0]     constant_24,
   input [31:0]     constant_25,
   input [31:0]     constant_26,
   input [31:0]     constant_27,
   input [31:0]     constant_28,
   input [31:0]     constant_29,
   input [31:0]     constant_30,
   input [31:0]     constant_31,
   input [31:0]     constant_32,
   input [31:0]     constant_33,
   input [31:0]     constant_34,
   input [31:0]     constant_35,
   input [31:0]     constant_36,
   input [31:0]     constant_37,
   input [31:0]     constant_38,
   input [31:0]     constant_39,
   input [31:0]     constant_40,
   input [31:0]     constant_41,
   input [31:0]     constant_42,
   input [31:0]     constant_43,
   input [31:0]     constant_44,
   input [31:0]     constant_45,
   input [31:0]     constant_46,
   input [31:0]     constant_47,
   input [31:0]     constant_48,
   input [31:0]     constant_49,
   input [31:0]     constant_50,
   input [31:0]     constant_51,
   input [31:0]     constant_52,
   input [31:0]     constant_53,
   input [31:0]     constant_54,
   input [31:0]     constant_55,
   input [31:0]     constant_56,
   input [31:0]     constant_57,
   input [31:0]     constant_58,
   input [31:0]     constant_59,
   input [31:0]     constant_60,
   input [31:0]     constant_61,
   input [31:0]     constant_62,
   input [31:0]     constant_63,
   input [31:0]     constant_64,
   input [31:0]     constant_65,
   input [31:0]     constant_66,
   input [31:0]     constant_67,
   input [31:0]     constant_68,
   input [31:0]     constant_69,
   input [31:0]     constant_70,
   input [31:0]     constant_71,
   input [31:0]     constant_72,
   input [31:0]     constant_73,
   input [31:0]     constant_74,
   input [31:0]     constant_75,
   input [31:0]     constant_76,
   input [31:0]     constant_77,
   input [31:0]     constant_78,
   input [31:0]     constant_79,
   input [31:0]     constant_80,
   input [31:0]     constant_81,
   input [31:0]     constant_82,
   input [31:0]     constant_83,
   input [31:0]     constant_84,
   input [31:0]     constant_85,
   input [31:0]     constant_86,
   input [31:0]     constant_87,
   input [31:0]     constant_88,
   input [31:0]     constant_89,
   input [31:0]     constant_90,
   input [31:0]     constant_91,
   input [31:0]     constant_92,
   input [31:0]     constant_93,
   input [31:0]     constant_94,
   input [31:0]     constant_95,
   input [31:0]                    delay0,
   input [31:0]                    delay1,
   input [31:0]                    delay2,
   input [31:0]                    delay3,
   input [31:0]                    delay4,
   input [31:0]                    delay5,
   input [31:0]                    delay6,
   input [31:0]                    delay7,
   input [31:0]                    delay8,
   input [31:0]                    delay9,
   input [31:0]                    delay10,
   input [31:0]                    delay11,
   input [31:0]                    delay12,
   input [31:0]                    delay13,
   input [31:0]                    delay14,
   input [31:0]                    delay15,
   input [31:0]                    delay16,
   input [31:0]                    delay17,
   input [31:0]                    delay18,
   input [31:0]                    delay19,
   input [31:0]                    delay20,
   input [31:0]                    delay21,
   input [31:0]                    delay22,
   input [31:0]                    delay23,
   input [31:0]                    delay24,
   input [31:0]                    delay25,
   input [31:0]                    delay26,
   input [31:0]                    delay27,
   input [31:0]                    delay28,
   input [31:0]                    delay29,
   input [31:0]                    delay30,
   input [31:0]                    delay31,
   input [31:0]                    delay32,
   input [31:0]                    delay33,
   input [31:0]                    delay34,
   input [31:0]                    delay35,
   input [31:0]                    delay36,
   input [31:0]                    delay37,
   input [31:0]                    delay38,
   input [31:0]                    delay39,
   input [31:0]                    delay40,
   input [31:0]                    delay41,
   input [31:0]                    delay42,
   input [31:0]                    delay43,
   input                           clk,
   input                           rst
   );

wire wor_ready;

wire [31:0] unitRdataFinal;
reg [31:0] stateRead;

// Memory access
wire [76:0] unitDone;

assign done = &unitDone;

wire [31:0] output_0_0 , output_1_0 , output_2_0 , output_3_0 , output_4_0 , output_5_0 , output_6_0 , output_7_0 , output_8_0 , output_9_0 , output_10_0 , output_11_0 , output_12_0 , output_13_0 , output_14_0 , output_15_0 , output_16_0 , output_17_0 , output_18_0 , output_19_0 , output_20_0 , output_21_0 , output_22_0 , output_23_0 , output_24_0 , output_25_0 , output_26_0 , output_27_0 , output_28_0 , output_29_0 , output_30_0 , output_31_0 , unused_32 , output_33_0 , output_34_0 , output_35_0 , output_36_0 , output_37_0 , output_38_0 , output_39_0 , output_40_0 , output_41_0 , output_42_0 , output_43_0 , output_44_0 , output_45_0 , output_46_0 , output_47_0 , output_48_0 , output_49_0 , output_50_0 , output_51_0 , output_52_0 , output_53_0 , output_54_0 , output_55_0 , output_56_0 , output_57_0 , output_58_0 , output_59_0 , output_60_0 , output_61_0 , output_62_0 , output_63_0 , output_64_0 , output_65_0 , output_66_0 , output_67_0 , output_68_0 , output_69_0 , output_70_0 , output_71_0 , output_72_0 , output_73_0 , output_74_0 , output_75_0 , output_76_0 ;

// Memory mapped
circuitInput circuitInput_0 (
      .in0(in0),
      .out0(output_0_0),
      .run(run),
      .done(unitDone[0]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_1 (
      .in0(in1),
      .out0(output_1_0),
      .run(run),
      .done(unitDone[1]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_2 (
      .in0(in2),
      .out0(output_2_0),
      .run(run),
      .done(unitDone[2]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_3 (
      .in0(in3),
      .out0(output_3_0),
      .run(run),
      .done(unitDone[3]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_4 (
      .in0(in4),
      .out0(output_4_0),
      .run(run),
      .done(unitDone[4]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_5 (
      .in0(in5),
      .out0(output_5_0),
      .run(run),
      .done(unitDone[5]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_6 (
      .in0(in6),
      .out0(output_6_0),
      .run(run),
      .done(unitDone[6]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_7 (
      .in0(in7),
      .out0(output_7_0),
      .run(run),
      .done(unitDone[7]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_8 (
      .in0(in8),
      .out0(output_8_0),
      .run(run),
      .done(unitDone[8]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_9 (
      .in0(in9),
      .out0(output_9_0),
      .run(run),
      .done(unitDone[9]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_10 (
      .in0(in10),
      .out0(output_10_0),
      .run(run),
      .done(unitDone[10]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_11 (
      .in0(in11),
      .out0(output_11_0),
      .run(run),
      .done(unitDone[11]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_12 (
      .in0(in12),
      .out0(output_12_0),
      .run(run),
      .done(unitDone[12]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_13 (
      .in0(in13),
      .out0(output_13_0),
      .run(run),
      .done(unitDone[13]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_14 (
      .in0(in14),
      .out0(output_14_0),
      .run(run),
      .done(unitDone[14]),
      .clk(clk),
      .rst(rst)
   );

circuitInput circuitInput_15 (
      .in0(in15),
      .out0(output_15_0),
      .run(run),
      .done(unitDone[15]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_16 (
      .out0(output_16_0),
      .in0(output_0_0),
      .in1(output_14_0),
      .in2(output_9_0),
      .in3(output_1_0),
      .constant_0(constant_0),
      .constant_1(constant_1),
      .constant_2(constant_2),
      .constant_3(constant_3),
      .constant_4(constant_4),
      .constant_5(constant_5),
      .run(run),
      .done(unitDone[16]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_17 (
      .out0(output_17_0),
      .in0(output_1_0),
      .in1(output_15_0),
      .in2(output_10_0),
      .in3(output_2_0),
      .constant_0(constant_6),
      .constant_1(constant_7),
      .constant_2(constant_8),
      .constant_3(constant_9),
      .constant_4(constant_10),
      .constant_5(constant_11),
      .run(run),
      .done(unitDone[17]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_18 (
      .out0(output_18_0),
      .in0(output_16_0),
      .in1(output_11_0),
      .in2(output_3_0),
      .in3(output_76_0),
      .constant_0(constant_12),
      .constant_1(constant_13),
      .constant_2(constant_14),
      .constant_3(constant_15),
      .constant_4(constant_16),
      .constant_5(constant_17),
      .run(run),
      .done(unitDone[18]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_19 (
      .out0(output_19_0),
      .in0(output_3_0),
      .in1(output_17_0),
      .in2(output_12_0),
      .in3(output_4_0),
      .constant_0(constant_18),
      .constant_1(constant_19),
      .constant_2(constant_20),
      .constant_3(constant_21),
      .constant_4(constant_22),
      .constant_5(constant_23),
      .run(run),
      .done(unitDone[19]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_20 (
      .out0(output_20_0),
      .in0(output_18_0),
      .in1(output_13_0),
      .in2(output_5_0),
      .in3(output_75_0),
      .constant_0(constant_24),
      .constant_1(constant_25),
      .constant_2(constant_26),
      .constant_3(constant_27),
      .constant_4(constant_28),
      .constant_5(constant_29),
      .run(run),
      .done(unitDone[20]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_21 (
      .out0(output_21_0),
      .in0(output_5_0),
      .in1(output_19_0),
      .in2(output_6_0),
      .in3(output_60_0),
      .constant_0(constant_30),
      .constant_1(constant_31),
      .constant_2(constant_32),
      .constant_3(constant_33),
      .constant_4(constant_34),
      .constant_5(constant_35),
      .run(run),
      .done(unitDone[21]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_22 (
      .out0(output_22_0),
      .in0(output_20_0),
      .in1(output_7_0),
      .in2(output_57_0),
      .in3(output_74_0),
      .constant_0(constant_36),
      .constant_1(constant_37),
      .constant_2(constant_38),
      .constant_3(constant_39),
      .constant_4(constant_40),
      .constant_5(constant_41),
      .run(run),
      .done(unitDone[22]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_23 (
      .out0(output_23_0),
      .in0(output_7_0),
      .in1(output_21_0),
      .in2(output_8_0),
      .in3(output_54_0),
      .constant_0(constant_42),
      .constant_1(constant_43),
      .constant_2(constant_44),
      .constant_3(constant_45),
      .constant_4(constant_46),
      .constant_5(constant_47),
      .run(run),
      .done(unitDone[23]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_24 (
      .out0(output_24_0),
      .in0(output_22_0),
      .in1(output_52_0),
      .in2(output_71_0),
      .in3(output_73_0),
      .constant_0(constant_48),
      .constant_1(constant_49),
      .constant_2(constant_50),
      .constant_3(constant_51),
      .constant_4(constant_52),
      .constant_5(constant_53),
      .run(run),
      .done(unitDone[24]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_25 (
      .out0(output_25_0),
      .in0(output_23_0),
      .in1(output_50_0),
      .in2(output_69_0),
      .in3(output_72_0),
      .constant_0(constant_54),
      .constant_1(constant_55),
      .constant_2(constant_56),
      .constant_3(constant_57),
      .constant_4(constant_58),
      .constant_5(constant_59),
      .run(run),
      .done(unitDone[25]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_26 (
      .out0(output_26_0),
      .in0(output_24_0),
      .in1(output_48_0),
      .in2(output_67_0),
      .in3(output_70_0),
      .constant_0(constant_60),
      .constant_1(constant_61),
      .constant_2(constant_62),
      .constant_3(constant_63),
      .constant_4(constant_64),
      .constant_5(constant_65),
      .run(run),
      .done(unitDone[26]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_27 (
      .out0(output_27_0),
      .in0(output_25_0),
      .in1(output_46_0),
      .in2(output_65_0),
      .in3(output_68_0),
      .constant_0(constant_66),
      .constant_1(constant_67),
      .constant_2(constant_68),
      .constant_3(constant_69),
      .constant_4(constant_70),
      .constant_5(constant_71),
      .run(run),
      .done(unitDone[27]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_28 (
      .out0(output_28_0),
      .in0(output_26_0),
      .in1(output_44_0),
      .in2(output_63_0),
      .in3(output_66_0),
      .constant_0(constant_72),
      .constant_1(constant_73),
      .constant_2(constant_74),
      .constant_3(constant_75),
      .constant_4(constant_76),
      .constant_5(constant_77),
      .run(run),
      .done(unitDone[28]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_29 (
      .out0(output_29_0),
      .in0(output_27_0),
      .in1(output_42_0),
      .in2(output_61_0),
      .in3(output_64_0),
      .constant_0(constant_78),
      .constant_1(constant_79),
      .constant_2(constant_80),
      .constant_3(constant_81),
      .constant_4(constant_82),
      .constant_5(constant_83),
      .run(run),
      .done(unitDone[29]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_30 (
      .out0(output_30_0),
      .in0(output_28_0),
      .in1(output_40_0),
      .in2(output_58_0),
      .in3(output_62_0),
      .constant_0(constant_84),
      .constant_1(constant_85),
      .constant_2(constant_86),
      .constant_3(constant_87),
      .constant_4(constant_88),
      .constant_5(constant_89),
      .run(run),
      .done(unitDone[30]),
      .clk(clk),
      .rst(rst)
   );

M_Stage M_Stage_31 (
      .out0(output_31_0),
      .in0(output_29_0),
      .in1(output_38_0),
      .in2(output_55_0),
      .in3(output_59_0),
      .constant_0(constant_90),
      .constant_1(constant_91),
      .constant_2(constant_92),
      .constant_3(constant_93),
      .constant_4(constant_94),
      .constant_5(constant_95),
      .run(run),
      .done(unitDone[31]),
      .clk(clk),
      .rst(rst)
   );

circuitOutput circuitOutput_32 (
      .out0(out0),
      .out1(out1),
      .out2(out2),
      .out3(out3),
      .out4(out4),
      .out5(out5),
      .out6(out6),
      .out7(out7),
      .out8(out8),
      .out9(out9),
      .out10(out10),
      .out11(out11),
      .out12(out12),
      .out13(out13),
      .out14(out14),
      .out15(out15),
      .in0(output_30_0),
      .in1(output_31_0),
      .in2(output_33_0),
      .in3(output_34_0),
      .in4(output_35_0),
      .in5(output_36_0),
      .in6(output_37_0),
      .in7(output_39_0),
      .in8(output_41_0),
      .in9(output_43_0),
      .in10(output_45_0),
      .in11(output_47_0),
      .in12(output_49_0),
      .in13(output_51_0),
      .in14(output_53_0),
      .in15(output_56_0),
      .run(run),
      .done(unitDone[32]),
      .clk(clk),
      .rst(rst)
   );

delay delay_33 (
      .out0(output_33_0),
      .in0(output_29_0),
      .delay0(delay0),
      .run(run),
      .done(unitDone[33]),
      .clk(clk),
      .rst(rst)
   );

delay delay_34 (
      .out0(output_34_0),
      .in0(output_28_0),
      .delay0(delay1),
      .run(run),
      .done(unitDone[34]),
      .clk(clk),
      .rst(rst)
   );

delay delay_35 (
      .out0(output_35_0),
      .in0(output_27_0),
      .delay0(delay2),
      .run(run),
      .done(unitDone[35]),
      .clk(clk),
      .rst(rst)
   );

delay delay_36 (
      .out0(output_36_0),
      .in0(output_26_0),
      .delay0(delay3),
      .run(run),
      .done(unitDone[36]),
      .clk(clk),
      .rst(rst)
   );

delay delay_37 (
      .out0(output_37_0),
      .in0(output_25_0),
      .delay0(delay4),
      .run(run),
      .done(unitDone[37]),
      .clk(clk),
      .rst(rst)
   );

delay delay_38 (
      .out0(output_38_0),
      .in0(output_24_0),
      .delay0(delay5),
      .run(run),
      .done(unitDone[38]),
      .clk(clk),
      .rst(rst)
   );

delay delay_39 (
      .out0(output_39_0),
      .in0(output_24_0),
      .delay0(delay6),
      .run(run),
      .done(unitDone[39]),
      .clk(clk),
      .rst(rst)
   );

delay delay_40 (
      .out0(output_40_0),
      .in0(output_23_0),
      .delay0(delay7),
      .run(run),
      .done(unitDone[40]),
      .clk(clk),
      .rst(rst)
   );

delay delay_41 (
      .out0(output_41_0),
      .in0(output_23_0),
      .delay0(delay8),
      .run(run),
      .done(unitDone[41]),
      .clk(clk),
      .rst(rst)
   );

delay delay_42 (
      .out0(output_42_0),
      .in0(output_22_0),
      .delay0(delay9),
      .run(run),
      .done(unitDone[42]),
      .clk(clk),
      .rst(rst)
   );

delay delay_43 (
      .out0(output_43_0),
      .in0(output_22_0),
      .delay0(delay10),
      .run(run),
      .done(unitDone[43]),
      .clk(clk),
      .rst(rst)
   );

delay delay_44 (
      .out0(output_44_0),
      .in0(output_21_0),
      .delay0(delay11),
      .run(run),
      .done(unitDone[44]),
      .clk(clk),
      .rst(rst)
   );

delay delay_45 (
      .out0(output_45_0),
      .in0(output_21_0),
      .delay0(delay12),
      .run(run),
      .done(unitDone[45]),
      .clk(clk),
      .rst(rst)
   );

delay delay_46 (
      .out0(output_46_0),
      .in0(output_20_0),
      .delay0(delay13),
      .run(run),
      .done(unitDone[46]),
      .clk(clk),
      .rst(rst)
   );

delay delay_47 (
      .out0(output_47_0),
      .in0(output_20_0),
      .delay0(delay14),
      .run(run),
      .done(unitDone[47]),
      .clk(clk),
      .rst(rst)
   );

delay delay_48 (
      .out0(output_48_0),
      .in0(output_19_0),
      .delay0(delay15),
      .run(run),
      .done(unitDone[48]),
      .clk(clk),
      .rst(rst)
   );

delay delay_49 (
      .out0(output_49_0),
      .in0(output_19_0),
      .delay0(delay16),
      .run(run),
      .done(unitDone[49]),
      .clk(clk),
      .rst(rst)
   );

delay delay_50 (
      .out0(output_50_0),
      .in0(output_18_0),
      .delay0(delay17),
      .run(run),
      .done(unitDone[50]),
      .clk(clk),
      .rst(rst)
   );

delay delay_51 (
      .out0(output_51_0),
      .in0(output_18_0),
      .delay0(delay18),
      .run(run),
      .done(unitDone[51]),
      .clk(clk),
      .rst(rst)
   );

delay delay_52 (
      .out0(output_52_0),
      .in0(output_17_0),
      .delay0(delay19),
      .run(run),
      .done(unitDone[52]),
      .clk(clk),
      .rst(rst)
   );

delay delay_53 (
      .out0(output_53_0),
      .in0(output_17_0),
      .delay0(delay20),
      .run(run),
      .done(unitDone[53]),
      .clk(clk),
      .rst(rst)
   );

delay delay_54 (
      .out0(output_54_0),
      .in0(output_16_0),
      .delay0(delay21),
      .run(run),
      .done(unitDone[54]),
      .clk(clk),
      .rst(rst)
   );

delay delay_55 (
      .out0(output_55_0),
      .in0(output_16_0),
      .delay0(delay22),
      .run(run),
      .done(unitDone[55]),
      .clk(clk),
      .rst(rst)
   );

delay delay_56 (
      .out0(output_56_0),
      .in0(output_16_0),
      .delay0(delay23),
      .run(run),
      .done(unitDone[56]),
      .clk(clk),
      .rst(rst)
   );

delay delay_57 (
      .out0(output_57_0),
      .in0(output_15_0),
      .delay0(delay24),
      .run(run),
      .done(unitDone[57]),
      .clk(clk),
      .rst(rst)
   );

delay delay_58 (
      .out0(output_58_0),
      .in0(output_15_0),
      .delay0(delay25),
      .run(run),
      .done(unitDone[58]),
      .clk(clk),
      .rst(rst)
   );

delay delay_59 (
      .out0(output_59_0),
      .in0(output_15_0),
      .delay0(delay26),
      .run(run),
      .done(unitDone[59]),
      .clk(clk),
      .rst(rst)
   );

delay delay_60 (
      .out0(output_60_0),
      .in0(output_14_0),
      .delay0(delay27),
      .run(run),
      .done(unitDone[60]),
      .clk(clk),
      .rst(rst)
   );

delay delay_61 (
      .out0(output_61_0),
      .in0(output_14_0),
      .delay0(delay28),
      .run(run),
      .done(unitDone[61]),
      .clk(clk),
      .rst(rst)
   );

delay delay_62 (
      .out0(output_62_0),
      .in0(output_14_0),
      .delay0(delay29),
      .run(run),
      .done(unitDone[62]),
      .clk(clk),
      .rst(rst)
   );

delay delay_63 (
      .out0(output_63_0),
      .in0(output_13_0),
      .delay0(delay30),
      .run(run),
      .done(unitDone[63]),
      .clk(clk),
      .rst(rst)
   );

delay delay_64 (
      .out0(output_64_0),
      .in0(output_13_0),
      .delay0(delay31),
      .run(run),
      .done(unitDone[64]),
      .clk(clk),
      .rst(rst)
   );

delay delay_65 (
      .out0(output_65_0),
      .in0(output_12_0),
      .delay0(delay32),
      .run(run),
      .done(unitDone[65]),
      .clk(clk),
      .rst(rst)
   );

delay delay_66 (
      .out0(output_66_0),
      .in0(output_12_0),
      .delay0(delay33),
      .run(run),
      .done(unitDone[66]),
      .clk(clk),
      .rst(rst)
   );

delay delay_67 (
      .out0(output_67_0),
      .in0(output_11_0),
      .delay0(delay34),
      .run(run),
      .done(unitDone[67]),
      .clk(clk),
      .rst(rst)
   );

delay delay_68 (
      .out0(output_68_0),
      .in0(output_11_0),
      .delay0(delay35),
      .run(run),
      .done(unitDone[68]),
      .clk(clk),
      .rst(rst)
   );

delay delay_69 (
      .out0(output_69_0),
      .in0(output_10_0),
      .delay0(delay36),
      .run(run),
      .done(unitDone[69]),
      .clk(clk),
      .rst(rst)
   );

delay delay_70 (
      .out0(output_70_0),
      .in0(output_10_0),
      .delay0(delay37),
      .run(run),
      .done(unitDone[70]),
      .clk(clk),
      .rst(rst)
   );

delay delay_71 (
      .out0(output_71_0),
      .in0(output_9_0),
      .delay0(delay38),
      .run(run),
      .done(unitDone[71]),
      .clk(clk),
      .rst(rst)
   );

delay delay_72 (
      .out0(output_72_0),
      .in0(output_9_0),
      .delay0(delay39),
      .run(run),
      .done(unitDone[72]),
      .clk(clk),
      .rst(rst)
   );

delay delay_73 (
      .out0(output_73_0),
      .in0(output_8_0),
      .delay0(delay40),
      .run(run),
      .done(unitDone[73]),
      .clk(clk),
      .rst(rst)
   );

delay delay_74 (
      .out0(output_74_0),
      .in0(output_6_0),
      .delay0(delay41),
      .run(run),
      .done(unitDone[74]),
      .clk(clk),
      .rst(rst)
   );

delay delay_75 (
      .out0(output_75_0),
      .in0(output_4_0),
      .delay0(delay42),
      .run(run),
      .done(unitDone[75]),
      .clk(clk),
      .rst(rst)
   );

delay delay_76 (
      .out0(output_76_0),
      .in0(output_2_0),
      .delay0(delay43),
      .run(run),
      .done(unitDone[76]),
      .clk(clk),
      .rst(rst)
   );

endmodule
